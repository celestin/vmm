class test extends vmm_test;

   function new(string name);
      super.new(name);
   endfunction

   // Lab 3 - Create the configure_test_ph() method
   // ToDo


endclass
test t_random = new("test");
