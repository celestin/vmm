James Chang                                           J a m e s   C h a n g                      J a m e s   C h a n g                                ��O    