program regfile_self_check;

endprogram: regfile_self_check