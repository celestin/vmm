`include "TR.sv"
`include "XACT.sv"
`include "MON.sv"
`include "SCBRD_CB.sv"
//`include "COV.sv"
`include "SB.sv"
