`include "test_cfg.sv"
`include "scoreboard.sv"
`include "coverage.sv"
`include "dut_env.sv"

