program test;

initial
begin
   top.env.run();
end
endprogram
